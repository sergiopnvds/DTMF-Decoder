LIBRARY ieee;
library std;
use std.textio.all;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
use ieee.std_logic_textio.all;

ENTITY tb_dtmf_top IS
END tb_dtmf_top;
 
ARCHITECTURE behavior OF tb_dtmf_top IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT dtmf_top
    PORT(
         clk : IN  std_logic;
         inputSignal : IN  signed(31 downto 0);
			outputTop : OUT  signed(6 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal inputSignal : signed(31 downto 0) := (others => '0');

 	--Outputs
   signal outputTop : signed(6 downto 0);

   -- Clock period definitions
   constant clk_period : time := 125 us;
	
	
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: dtmf_top PORT MAP (
          clk => clk,
          outputTop => outputTop,
          inputSignal => inputSignal
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   -- Stimulus process
   stim_proc: process

	file fichero_seno : text open read_mode is "C:\Users\Abinarios.txt"; 
	variable linea : line;
	variable valor : std_logic_vector(31 downto 0);
	
   begin		
		--if(clk ' event and clk = '1') then
		  wait for clk_period/2;
		  while not(endfile(fichero_seno)) loop
		    readline(fichero_seno, linea);
			 read(linea, valor);
			 inputSignal <= signed(valor);
			 wait for clk_period;
		  end loop;
		--end if;

--begin	
--	wait for 100ns;
--inputSignal<="00000000000000001010100100000100"; wait for 125 us;
--inputSignal<="00000000000000011010010101110000";wait for 125 us;
--inputSignal<="00000000000000010011101111010101";wait for 125 us;
--
--inputSignal<="11111111111111111000110101100110";wait for 125 us;
--
--inputSignal<="11111111111111100110011100011100";wait for 125 us;
--
--inputSignal<="11111111111111101101101100111000";wait for 125 us;
--
--inputSignal<="11111111111111111110001110011110";wait for 125 us;
--
--inputSignal<="11111111111111111111010100010110";wait for 125 us;
--
--inputSignal<="11111111111111110011100111101001";wait for 125 us;
--
--inputSignal<="11111111111111110100000110110100";wait for 125 us;
--
--inputSignal<="00000000000000001001111011011111";wait for 125 us;
--
--inputSignal<="00000000000000011110011100000000";wait for 125 us;
--
--inputSignal<="00000000000000011001000101111010";wait for 125 us;
--
--inputSignal<="00000000000000000001001011110110";wait for 125 us;
--
--inputSignal<="11111111111111110011100000011001";wait for 125 us;
--
--inputSignal<="11111111111111111010101101111111";wait for 125 us;
--
--inputSignal<="00000000000000000010101100111001";wait for 125 us;
--
--inputSignal<="11111111111111111000001101110100";wait for 125 us;
--
--inputSignal<="11111111111111100110101110100000";wait for 125 us;
--
--inputSignal<="11111111111111101001000001110100";wait for 125 us;
--
--inputSignal<="00000000000000000010010111111100";wait for 125 us;
--
--inputSignal<="00000000000000010111111010000001";wait for 125 us;
--
--inputSignal<="00000000000000010100010110010000";wait for 125 us;
--
--inputSignal<="00000000000000000011101010110011";wait for 125 us;
--
--inputSignal<="11111111111111111111111100011010";wait for 125 us;
--
--inputSignal<="00000000000000001011011000011111";wait for 125 us;
--
--inputSignal<="00000000000000001110000101001001";wait for 125 us;
--
--inputSignal<="11111111111111111010011100000001";wait for 125 us;
--
--inputSignal<="11111111111111100011011110010000";wait for 125 us;
--
--inputSignal<="11111111111111100100010000100001";wait for 125 us;
--
--inputSignal<="11111111111111111010110111001001";wait for 125 us;
--
--inputSignal<="00000000000000001011010110010100";wait for 125 us;
--
--inputSignal<="00000000000000000110011110100101";wait for 125 us;
--
--inputSignal<="11111111111111111101000100110010";wait for 125 us;
--
--inputSignal<="00000000000000000101000100010100";wait for 125 us;
--
--inputSignal<="00000000000000010111100111110100";wait for 125 us;
--
--inputSignal<="00000000000000011001100101000100";wait for 125 us;
--
--inputSignal<="00000000000000000010100000010111";wait for 125 us;
--
--inputSignal<="11111111111111101010011010011111";wait for 125 us;
--
--inputSignal<="11111111111111101010000001011100";wait for 125 us;
--
--inputSignal<="11111111111111111010001110100111";wait for 125 us;
--
--inputSignal<="00000000000000000000100000110111";wait for 125 us;
--
--inputSignal<="11111111111111110101111000000010";wait for 125 us;
--
--inputSignal<="11111111111111110000010001001001";wait for 125 us;
--
--inputSignal<="00000000000000000001001101010111";wait for 125 us;
--
--inputSignal<="00000000000000011001111011100101";wait for 125 us;
--
--inputSignal<="00000000000000011101101111111001";wait for 125 us;
--
--inputSignal<="00000000000000001001001010010001";wait for 125 us;
--
--inputSignal<="11111111111111110110010010100011";wait for 125 us;
--
--inputSignal<="11111111111111111000011101110100";wait for 125 us;
--
--inputSignal<="00000000000000000010110011010100";wait for 125 us;
--
--inputSignal<="11111111111111111101011111111000";wait for 125 us;
--
--inputSignal<="11111111111111101010100010100101";wait for 125 us;
--
--inputSignal<="11111111111111100100011111110111";wait for 125 us;
--
--inputSignal<="11111111111111111000101001111011";wait for 125 us;
--
--inputSignal<="00000000000000010010101001000001";wait for 125 us;
--
--inputSignal<="00000000000000010111000111000101";wait for 125 us;
--
--inputSignal<="00000000000000001000000000100010";wait for 125 us;
--
--inputSignal<="11111111111111111111010110001101";wait for 125 us;
--
--inputSignal<="00000000000000001000101011111001";wait for 125 us;
--
--inputSignal<="00000000000000010000110101001010";wait for 125 us;
--
--inputSignal<="00000000000000000011000000101101";wait for 125 us;
--
--inputSignal<="11111111111111101001010001101100";wait for 125 us;
--
--inputSignal<="11111111111111100000111101000100";wait for 125 us;
--
--inputSignal<="11111111111111110010110111010111";wait for 125 us;
--
--inputSignal<="00000000000000000111100110010011";wait for 125 us;
--
--inputSignal<="00000000000000001000010111111110";wait for 125 us;
--
--inputSignal<="11111111111111111101101000101010";wait for 125 us;
--
--inputSignal<="00000000000000000000001010110000";wait for 125 us;
--
--inputSignal<="00000000000000010010110111110111";wait for 125 us;
--
--inputSignal<="00000000000000011100101100111110";wait for 125 us;
--
--inputSignal<="00000000000000001100000000110101";wait for 125 us;
--
--inputSignal<="11111111111111110000110111010010";wait for 125 us;
--
--inputSignal<="11111111111111101000010100010111";wait for 125 us;
--
--inputSignal<="11111111111111110101101101000111";wait for 125 us;
--
--inputSignal<="00000000000000000000011101000100";wait for 125 us;
--
--inputSignal<="11111111111111111000110110011010";wait for 125 us;
--
--inputSignal<="11111111111111101110100111110111";wait for 125 us;
--
--inputSignal<="11111111111111111001000000111111";wait for 125 us;
--
--inputSignal<="00000000000000010010111111110111";wait for 125 us;
--
--inputSignal<="00000000000000011111100101110000";wait for 125 us;
--
--inputSignal<="00000000000000010000111100011011";wait for 125 us;
--
--inputSignal<="11111111111111111010111100101100";wait for 125 us;
--
--inputSignal<="11111111111111110111000100100001";wait for 125 us;
--
--inputSignal<="00000000000000000001101010010111";wait for 125 us;
--
--inputSignal<="00000000000000000001110111100100";wait for 125 us;
--
--inputSignal<="11111111111111110000000010101010";wait for 125 us;
--
--inputSignal<="11111111111111100010110101011110";wait for 125 us;
--
--inputSignal<="11111111111111101111100111011101";wait for 125 us;
--
--inputSignal<="00000000000000001011001010000010";wait for 125 us;
--
--inputSignal<="00000000000000010111101001000111";wait for 125 us;
--
--inputSignal<="00000000000000001100100010101011";wait for 125 us;
--
--inputSignal<="00000000000000000000000101101010";wait for 125 us;
--
--inputSignal<="00000000000000000101100110011101";wait for 125 us;
--
--inputSignal<="00000000000000010001011001000110";wait for 125 us;
--
--inputSignal<="00000000000000001010100110111111";wait for 125 us;
--
--inputSignal<="11111111111111110001001000111101";wait for 125 us;
--
--inputSignal<="11111111111111100000101001001011";wait for 125 us;
--
--inputSignal<="11111111111111101011100001111001";wait for 125 us;
--
--inputSignal<="00000000000000000010001000000100";wait for 125 us;
--
--inputSignal<="00000000000000001001001000111011";wait for 125 us;
--
--inputSignal<="11111111111111111111001111110111";wait for 125 us;
--
--inputSignal<="11111111111111111100011100100000";wait for 125 us;
--
--inputSignal<="00000000000000001100110100100011";wait for 125 us;
--
--inputSignal<="00000000000000011100111001001011";wait for 125 us;
--
--inputSignal<="00000000000000010100010101101111";wait for 125 us;
--
--inputSignal<="11111111111111111001001100101011";wait for 125 us;
--
--inputSignal<="11111111111111101001000010011011";wait for 125 us;
--
--inputSignal<="11111111111111110001010110000110";wait for 125 us;
--
--inputSignal<="11111111111111111111000010011000";wait for 125 us;
--
--inputSignal<="11111111111111111011111000010110";wait for 125 us;
--
--inputSignal<="11111111111111101111000101100101";wait for 125 us;
--
--inputSignal<="11111111111111110010001101000010";wait for 125 us;
--
--inputSignal<="00000000000000001010011011011001";wait for 125 us;
--
--inputSignal<="00000000000000011110010110001001";wait for 125 us;
--
--inputSignal<="00000000000000010111100110101000";wait for 125 us;
--
--inputSignal<="00000000000000000001000110110100";wait for 125 us;
--
--inputSignal<="11111111111111110111000010101110";wait for 125 us;
--
--inputSignal<="11111111111111111111101101001000";wait for 125 us;
--
--inputSignal<="00000000000000000100110110110000";wait for 125 us;
--
--inputSignal<="11111111111111110110011011101101";wait for 125 us;
--
--inputSignal<="11111111111111100100000101010101";wait for 125 us;
--
--inputSignal<="11111111111111101000001110010111";wait for 125 us;
--
--inputSignal<="00000000000000000010001011110111";wait for 125 us;
--
--inputSignal<="00000000000000010101101000011000";wait for 125 us;
--
--inputSignal<="00000000000000010000100010101011";wait for 125 us;
--
--inputSignal<="00000000000000000010001001000000";wait for 125 us;
--
--inputSignal<="00000000000000000010110001111111";wait for 125 us;
--
--inputSignal<="00000000000000001111111111100100";wait for 125 us;
--
--inputSignal<="00000000000000010000011110010100";wait for 125 us;
--
--inputSignal<="11111111111111111010001011001001";wait for 125 us;
--
--inputSignal<="11111111111111100011011010111010";wait for 125 us;
--
--inputSignal<="11111111111111100101110000100101";wait for 125 us;
--
--inputSignal<="11111111111111111011011100001100";wait for 125 us;
--
--inputSignal<="00000000000000001000010110100000";wait for 125 us;
--
--inputSignal<="00000000000000000001011001111010";wait for 125 us;
--
--inputSignal<="11111111111111111010001111111000";wait for 125 us;
--
--inputSignal<="00000000000000000110010011011001";wait for 125 us;
--
--inputSignal<="00000000000000011010010010000111";wait for 125 us;
--
--inputSignal<="00000000000000011010100110100100";wait for 125 us;
--
--inputSignal<="00000000000000000010100100100001";wait for 125 us;
--
--inputSignal<="11111111111111101100010101110110";wait for 125 us;
--
--inputSignal<="11111111111111101101111000101111";wait for 125 us;
--
--inputSignal<="11111111111111111100011010111110";wait for 125 us;
--
--inputSignal<="11111111111111111110010110010101";wait for 125 us;
--
--inputSignal<="11111111111111110001010011001110";wait for 125 us;
--
--inputSignal<="11111111111111101101011010011011";wait for 125 us;
--
--inputSignal<="00000000000000000001001011101001";wait for 125 us;
--inputSignal<="00000000000000011010000110100001";wait for 125 us;
--inputSignal<="00000000000000011100010010110011";wait for 125 us;
--inputSignal<="00000000000000001000001000101011";wait for 125 us;
--inputSignal<="11111111111111111000101100011010";wait for 125 us;
--inputSignal<="11111111111111111101100000000110";wait for 125 us;
--inputSignal<="00000000000000000110001111100101";wait for 125 us;
--inputSignal<="11111111111111111100110111100110";wait for 125 us;
--inputSignal<="11111111111111100111111100010010";wait for 125 us;
--inputSignal<="11111111111111100011010000000100";wait for 125 us;
--inputSignal<="11111111111111111000101010011000";wait for 125 us;
--inputSignal<="00000000000000010001000100111001";wait for 125 us;
--inputSignal<="00000000000000010011010010011101";wait for 125 us;
--inputSignal<="00000000000000000101001110000000";wait for 125 us;
--inputSignal<="00000000000000000000110010001100";wait for 125 us;
--inputSignal<="00000000000000001101000111000001";wait for 125 us;
--inputSignal<="00000000000000010100000110100010";wait for 125 us;
--inputSignal<="00000000000000000011011000000111";wait for 125 us;
--inputSignal<="11111111111111101001000001011010";wait for 125 us;
--inputSignal<="11111111111111100010010011111100";wait for 125 us;
--inputSignal<="11111111111111110100010001011000";wait for 125 us;
--inputSignal<="00000000000000000101110100101001";wait for 125 us;
--inputSignal<="00000000000000000011011111110111";wait for 125 us;
--inputSignal<="11111111111111111001101001111001";wait for 125 us;
--inputSignal<="00000000000000000000001001010111";wait for 125 us;
--inputSignal<="00000000000000010101010100110011";wait for 125 us;
--inputSignal<="00000000000000011110001010100000";wait for 125 us;
--inputSignal<="00000000000000001011111111000111";wait for 125 us;
--inputSignal<="11111111111111110010000100000111";wait for 125 us;
--inputSignal<="11111111111111101100000000010100";wait for 125 us;
--inputSignal<="11111111111111111001000000100000";wait for 125 us;
--inputSignal<="11111111111111111111110001111000";wait for 125 us;
--inputSignal<="11111111111111110100101100010100";wait for 125 us;
--inputSignal<="11111111111111101010111111101110";wait for 125 us;
--inputSignal<="11111111111111111000010001011010";wait for 125 us;
--inputSignal<="00000000000000010011010010101101";wait for 125 us;
--inputSignal<="00000000000000011110010111101100";wait for 125 us;
--inputSignal<="00000000000000001111001110100101";wait for 125 us;
--inputSignal<="11111111111111111100000101000011";wait for 125 us;
--inputSignal<="11111111111111111011101011000001";wait for 125 us;
--inputSignal<="00000000000000000110000101110010";wait for 125 us;
--inputSignal<="00000000000000000010100100010110";wait for 125 us;
--inputSignal<="11111111111111101101110100100010";wait for 125 us;
--inputSignal<="11111111111111100001001011101000";wait for 125 us;
--inputSignal<="11111111111111101111100111001101";wait for 125 us;
--inputSignal<="00000000000000001010010011101011";wait for 125 us;
--inputSignal<="00000000000000010100001011010010";wait for 125 us;
--inputSignal<="00000000000000001000110100100001";wait for 125 us;
--inputSignal<="11111111111111111111111111000110";wait for 125 us;
--inputSignal<="00000000000000001001011000011101";wait for 125 us;
--inputSignal<="00000000000000010101010011001101";wait for 125 us;
--inputSignal<="00000000000000001011110000100011";wait for 125 us;
--inputSignal<="11111111111111110000110110110000";wait for 125 us;
--inputSignal<="11111111111111100001101100100011";wait for 125 us;
--inputSignal<="11111111111111101101011110101001";wait for 125 us;
--inputSignal<="00000000000000000001101000111000";wait for 125 us;
--inputSignal<="00000000000000000100111010111000";wait for 125 us;
--inputSignal<="11111111111111111010011110011011";wait for 125 us;
--inputSignal<="11111111111111111011000011110000";wait for 125 us;
--inputSignal<="00000000000000001110101110011111";wait for 125 us;
--inputSignal<="00000000000000011110101101001010";wait for 125 us;
--inputSignal<="00000000000000010100011010111010";wait for 125 us;
--inputSignal<="11111111111111111001101110001100";wait for 125 us;
--inputSignal<="11111111111111101100001101011010";wait for 125 us;
--inputSignal<="11111111111111110101011000010111";wait for 125 us;
--inputSignal<="11111111111111111111111010010111";wait for 125 us;
--11111111111111111000100100111110";wait for 125 us;
--11111111111111101010111111000100";wait for 125 us;
--11111111111111110000101000100110";wait for 125 us;
--00000000000000001010101001100010";wait for 125 us;
--00000000000000011101011110100100";wait for 125 us;
--00000000000000010101011111111111";wait for 125 us;
--00000000000000000000111110000101";wait for 125 us;
--11111111111111111010110010001100";wait for 125 us;
--00000000000000000100101101010001";wait for 125 us;
--00000000000000000110111010110100";wait for 125 us;
--11111111111111110100111011000001";wait for 125 us;
--11111111111111100010001010001010";wait for 125 us;
--11111111111111101000000001101110";wait for 125 us;
--00000000000000000001111100110111";wait for 125 us;
--00000000000000010010110100000110";wait for 125 us;
--00000000000000001100010011010010";wait for 125 us;
--00000000000000000000100001010101";wait for 125 us;
--00000000000000000101100000111010";wait for 125 us;
--00000000000000010100001100010001";wait for 125 us;
--00000000000000010010011101101011";wait for 125 us;
--11111111111111111010000100100111";wait for 125 us;
--11111111111111100100000110011000";wait for 125 us;
--11111111111111100111111100001010";wait for 125 us;
--11111111111111111100001010100000";wait for 125 us;
--00000000000000000101001010110001";wait for 125 us;
--11111111111111111100010010110011";wait for 125 us;
--11111111111111110111100010011000";wait for 125 us;
--00000000000000000111010110010001";wait for 125 us;
--00000000000000011100010000110111";wait for 125 us;
--00000000000000011010111100101001";wait for 125 us;
--00000000000000000010100011111001";wait for 125 us;
--11111111111111101110110000100000";wait for 125 us;
--11111111111111110010001110001000";wait for 125 us;
--11111111111111111110101111011011";wait for 125 us;
--11111111111111111100010000110011";wait for 125 us;
--11111111111111101101000111000001";wait for 125 us;
--11111111111111101011000001001000";wait for 125 us;
--00000000000000000001000111001000";wait for 125 us;
--00000000000000011001100110101011";wait for 125 us;
--00000000000000011010000111000001";wait for 125 us;
--00000000000000000110111000000101";wait for 125 us;
--11111111111111111011010000010100";wait for 125 us;
--00000000000000000010100110001110";wait for 125 us;
--00000000000000001001100011011001";wait for 125 us;
--11111111111111111100010110011110";wait for 125 us;
--11111111111111100101111110000101";wait for 125 us;
--11111111111111100010101111001110";wait for 125 us;
--11111111111111111000110111010110";wait for 125 us;
--00000000000000001111000101110100";wait for 125 us;
--00000000000000001110111110001000";wait for 125 us;
--00000000000000000010010000111010";wait for 125 us;
--00000000000000000010001010011101";wait for 125 us;
--00000000000000010001001011110011";wait for 125 us;
--00000000000000010110110111110101";wait for 125 us;
--00000000000000000011101010111010";wait for 125 us;
--11111111111111101001010110110101";wait for 125 us;
--11111111111111100100011011101010";wait for 125 us;
--11111111111111110110000000000111";wait for 125 us;
--00000000000000000011111011100010
--11111111111111111110100010101010
--11111111111111110101110100000001
--00000000000000000000000101101010
--00000000000000010111001101111001
--00000000000000011110110110101100
--00000000000000001011101001011000
--11111111111111110011100110101100
--11111111111111110000001100110100
--11111111111111111100100001000110
--11111111111111111111001001100110
--11111111111111110000110101111101
--11111111111111100111111001010110
--11111111111111110111101101100000
--00000000000000010011000101110011
--00000000000000011100010111110011
--00000000000000001101000110011110
--11111111111111111101010001101100
--00000000000000000000010111100111
--00000000000000001010011000011101
--00000000000000000011001111000010
--11111111111111101100000101010100
--11111111111111100000010100010000
--11111111111111110000000010000101
--00000000000000001001001101100001
--00000000000000010000001100111010
--00000000000000000100110110011101
--11111111111111111111110101111111
--00000000000000001100111001100101
--00000000000000011000101010110100
--00000000000000001100100111110100
--11111111111111110000111101100100
--11111111111111100011100001100001
--11111111111111101111111010110110
--00000000000000000001001001001100
--00000000000000000000100110000111
--11111111111111110101110101001010
--11111111111111111001110001000001
--00000000000000010000001110111111
--00000000000000011111101110110000
--00000000000000010011111110011011
--11111111111111111010011000111011
--11111111111111101111111000000100
--11111111111111111001101101001010
--00000000000000000000110100111111
--11111111111111110101011111100100
--11111111111111100111011010110111
--11111111111111101111011100010110
--00000000000000001010100101111011
--00000000000000011011110110110101
--00000000000000010010110101001111
--00000000000000000000110001100111
--11111111111111111110101000100101
--00000000000000001001100110001101
--00000000000000001000110101100011
--11111111111111110011101101111101
--11111111111111100001000000000110
--11111111111111101000011100100000
--00000000000000000001101011101100
--00000000000000001111100001111101
--00000000000000000111101110111100
--11111111111111111110110110011000
--00000000000000001000000100110000
--00000000000000010111110111101100
--00000000000000010011111111101100
--11111111111111111010001000001011
--11111111111111100101011111011000
--11111111111111101010101111110011
--11111111111111111101000001001010
--00000000000000000001111000011100
--11111111111111110111010001101000
--11111111111111110101000000111010
--00000000000000001000001011011110
--00000000000000011101100000111101
--00000000000000011010100110011111
--00000000000000000010011110000110
--11111111111111110001100110010001
--11111111111111110110111010100001
--00000000000000000001001000001011
--11111111111111111010010011101001
--11111111111111101001011010010000
--11111111111111101001001001011001
--00000000000000000001000000010011
--00000000000000011000011101000111
--00000000000000010111010000000000
--00000000000000000101011010010100
--11111111111111111101111001111001
--00000000000000000111100111110110
--00000000000000001100101001001101
--11111111111111111011111101000011
--11111111111111100100101011000011
--11111111111111100010111110011000
--11111111111111111001010000110111
--00000000000000001100101111010010
--00000000000000001010010001001101
--11111111111111111111001110000100
--00000000000000000011011100110001
--00000000000000010100110011101000
--00000000000000011001000100010101
--00000000000000000011111000010000
--11111111111111101010010001001010
--11111111111111100111010000110001
--11111111111111111000000000111111
--00000000000000000001111110001110
--11111111111111111001101000011111
--11111111111111110010001101011010
--00000000000000000000000000000000
--00000000000000011000100000010010
--00000000000000011110110000010100
--00000000000000001010111111110010
--11111111111111110101011100001101
--11111111111111110100110010111011
--00000000000000000000001001001010
--11111111111111111110100101001100
--11111111111111101101011001100010
--11111111111111100101011001111101
--11111111111111110111010110100100
--00000000000000010010011001110100
--00000000000000011001101001011010
--00000000000000001010100111010111
--11111111111111111110100000011101
--00000000000000000101000010100110
--00000000000000001110011011010000
--00000000000000000011110110010001
--11111111111111101010110111100100
--11111111111111100000010000110101
--11111111111111110000110111110001
--00000000000000000111111001101101
--00000000000000001011110100100100
--00000000000000000000101110111110
--11111111111111111111101010100110
--00000000000000010000000100001010
--00000000000000011011011010010101
--00000000000000001101001011000100
--11111111111111110001011100111000
--11111111111111100110000101000000
--11111111111111110010110010101100
--00000000000000000000101001111111
--11111111111111111100010001110000
--11111111111111110001011011101111
--11111111111111111000100110101010
--00000000000000010001010011111000
--00000000000000011111111100010001
--00000000000000010011000000101100
--11111111111111111011001011011010
--11111111111111110011111100010010
--11111111111111111110001101011011
--00000000000000000001110000110001
--11111111111111110010101101000010
--11111111111111100100011110110111
--11111111111111101110101010100101
--00000000000000001010010001000010
--00000000000000011001100001101110
--00000000000000001111101010100101
--00000000000000000000100001100010
--00000000000000000010011111100001
--00000000000000001110001111111010
--00000000000000001010100011100100
--11111111111111110010110110001100
--11111111111111100000101000111101
--11111111111111101001011110010001
--00000000000000000001011001001011
--00000000000000001011110111011111
--00000000000000000010111101001001
--11111111111111111101001010111001
--00000000000000001010011001011100
--00000000000000011010111011110110
--00000000000000010101000001100101
--11111111111111111010010101010110
--11111111111111100111100011011011
--11111111111111101110000111000100
--11111111111111111101111110111101
--11111111111111111110100101000000
--11111111111111110010011110101001
--11111111111111110010101111110001
--00000000000000001000110001111110
--00000000000000011110000000011101
--00000000000000011001100100011101
--00000000000000000010010010111100
--11111111111111110100110010010001
--11111111111111111011110110001110
--00000000000000000011100001010111
--11111111111111111000100001111011
--11111111111111100110010010111100
--11111111111111100111110110100001
--00000000000000000000110111110001
--00000000000000010110101011111011
--00000000000000010011110010011000
--00000000000000000011110001100011
--00000000000000000000100100101111
--00000000000000001100011100101100
--00000000000000001111011011110011
--11111111111111111011101011101101
--11111111111111100100000101000111
--11111111111111100011111101010010
--11111111111111111001110110101001
--00000000000000001010000101011010
--00000000000000000101010011011001
--11111111111111111100001010011100
--00000000000000000100100111001011
--00000000000000010111111000101000
--00000000000000011010101000010000
--00000000000000000011111111011000
--11111111111111101011101110100100
--11111111111111101010101110101011
--11111111111111111010010000111000
--00000000000000000000000000000000
--11111111111111110100111001011001
--11111111111111101110111100000110
--11111111111111111111111000110101
--00000000000000011001001010000100
--00000000000000011101110111011010
--00000000000000001010000011000110
--11111111111111110111100001011000
--11111111111111111001101011000101
--00000000000000000011110010110100
--11111111111111111110000101011110
--11111111111111101010011100100110
--11111111111111100011100101110001
--11111111111111110111001101100110
--00000000000000010001010000001100
--00000000000000010110010000111101
--00000000000000000111110101001001
--11111111111111111111101111001110
--00000000000000001001100100010011
--00000000000000010010000111011100
--00000000000000000100011000101111
--11111111111111101010001101000010
--11111111111111100001000001011111
--11111111111111110010000111001101
--00000000000000000110011010101001
--00000000000000000111001001100000
--11111111111111111100100100110010
--11111111111111111111011101010110
--00000000000000010010110011001001
--00000000000000011101011101001001
--00000000000000001101011000111111
--11111111111111110010010011100001
--11111111111111101001010010110010
--11111111111111110110000001101010
--00000000000000000000001100001101
--11111111111111111000000100110101
--11111111111111101101011001011100
--11111111111111110111100110110111
--00000000000000010001111011101100
--00000000000000011111010101011001
--00000000000000010001100011000000
--11111111111111111100000100000011
--11111111111111111000010011010001
--00000000000000000010110001110010
--00000000000000000010101100000100
--11111111111111110000010001110101
--11111111111111100010001111111001
--11111111111111101110010100111010
--00000000000000001001101011110100
--00000000000000010110100011001100
--00000000000000001100000101000100
--00000000000000000000001110001000
--00000000000000000110010000101101
--00000000000000010010100010101010
--00000000000000001100000001110011
--11111111111111110010010100110100
--11111111111111100001000101010001
--11111111111111101011000101100110
--00000000000000000001000110000101
--00000000000000000111111010110111
--11111111111111111110000101101101
--11111111111111111011100001101110
--00000000000000001100011011010110
--00000000000000011101010011101101
--00000000000000010101100001010110
--11111111111111111010101011011001
--11111111111111101010001110111110
--11111111111111110001111100100010
--11111111111111111111000010011101
--11111111111111111011010101110101
--11111111111111101110000001110000
--11111111111111110000110010111010
--00000000000000001001001001000111
--00000000000000011101101110101110
--00000000000000010111111000000001
--00000000000000000010000010010111
--11111111111111111000001111001000
--00000000000000000000111001001001
--00000000000000000101110110111110
--11111111111111110110111110011001
--11111111111111100011110110001000
--11111111111111100111001010111001
--00000000000000000000101110001010
--00000000000000010100010110001111
--00000000000000001111110011101111
--00000000000000000010000000010101
--00000000000000000011001100011100
--00000000000000010000111100110111
--00000000000000010001110110011010
--11111111111111111011100010011111
--11111111111111100100001101000100
--11111111111111100101101010011111
--11111111111111111010101000000011
--00000000000000000111001100101110
--00000000000000000000001100110111
--11111111111111111001001011000101
--00000000000000000101100111111010
--00000000000000011010010101111001
--00000000000000011011100000110101
--00000000000000000011111111101101
--11111111111111101101101100011011
--11111111111111101110101111101110
--11111111111111111100101100010000
--11111111111111111110000100001010
--11111111111111110000011101001001
--11111111111111101100000101101001
--11111111111111111111110000101011
--00000000000000011001001010011011
--00000000000000011100001101010101
--00000000000000001000110100100000
--11111111111111111001110010100101
--11111111111111111110101101010001
--00000000000000000111011000000001
--11111111111111111101101011000110
--11111111111111101000000011110100
--11111111111111100010011111111010
--11111111111111110111010011001100
--00000000000000001111101011001000
--00000000000000010010010100000000
--00000000000000000100110100001111
--00000000000000000000111011111010
--00000000000000001101110101010100
--00000000000000010101010110110110
--00000000000000000100110101010000
--11111111111111101010000110100000
--11111111111111100010100101000001
--11111111111111110011101110101010
--00000000000000000100110011000011
--00000000000000000010010011011100
--11111111111111111000011110101111
--11111111111111111111001110101111
--00000000000000010101000010001110
--00000000000000011110101111110100
--00000000000000001101010000111000
--11111111111111110011011111101111
--11111111111111101101000101100000
--11111111111111111001100010100011
--11111111111111111111110000101010
--11111111111111110100000110001111
--11111111111111101001110100111111
--11111111111111110110110011100101
--00000000000000010010000101101111
--00000000000000011101111011001001
--00000000000000001111100111011111
--11111111111111111101000001001001
--11111111111111111100110101110011
--00000000000000000111010010101111
--00000000000000000011100101001101
--11111111111111101110010001101100
--11111111111111100000110001101011
--11111111111111101110011100001101
--00000000000000001000110111100100
--00000000000000010011000000001101
--00000000000000001000001010011110
--11111111111111111111110111110101
--00000000000000001001110101111111
--00000000000000010110010111011010
--00000000000000001101001101100100
--11111111111111110010001010010110
--11111111111111100010010100001101
--11111111111111101101010000000101
--00000000000000000000110011001101
--00000000000000000011110010100111
--11111111111111111001010000100110
--11111111111111111001111101101100
--00000000000000001110000111010111
--00000000000000011110111011011010
--00000000000000010101011101111000
--11111111111111111011001001010110
--11111111111111101101011101011101
--11111111111111110110001010000000
--00000000000000000000001001111111

   end process;

END;

